`timescale 10ps / 1ps
module list_1(input input_tmp, output output_tmp);

exercise4tb e4tb ();
exercise5tb e5tb ();
exercise6tb e6tb ();
exercise7tb e7tb ();

endmodule 